module new #(
    parameters
) (
    ports
);
    
endmodule